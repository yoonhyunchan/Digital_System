module mux();


input IN1;
input IN2;


endmodule