module MEM();





endmodule