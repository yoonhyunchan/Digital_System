module ALU(ALUIN1, ALUIN2, ALUC, ALU_OUT);
    input [31:0] ALU_IN1;
    input [31:0] ALU_IN2;
    input ALUC;
    output reg [31:0] CLU_OUT;


    always @(posedge ALUC) begin
    end
    
endmodule