module tb();



endmodule