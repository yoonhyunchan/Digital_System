module SingleCpu(CLK);
    input CLK;



Vr_data_mem Vr_data_mem1(CLK, ADDR, RW, WD, RD);







endmodule