module IF_ID(Data, RST);

always @(Data or RST) begin
    
end



endmodule