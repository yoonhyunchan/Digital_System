module IF_ID(Data, RST);

    input Data;
    input RST;
    output reg Q;

always @(Data or RST) begin
    
end



endmodule