module MEM();


endmodule