module EX_MEM ();
    input nPC_M;




    
endmodule