module EX_MEM ();
    output reg nPC_M;
    output reg AOUT_M;
    output reg B_M;



    
endmodule