module IF_ID(Data, RST);

    input Data;
    input RST;

always @(Data or RST) begin
    
end



endmodule