module ALU(ALU_CIN, ALUIN1, ALUIN2, ALUC, ALU_OUT);
    input ALU_CIN;
    output reg CLU_OUT;
    

    // always @(*) begin
    // end
    
endmodule