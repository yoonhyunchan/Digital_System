module Control();




endmodule