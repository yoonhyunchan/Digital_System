module ID_EX();


    input RD1;
    input RD2;
    input signout;
    


endmodule