module MEM_WB ();
    
    output reg [31:0] MDR_W;
    output reg [31:0] AOUT_W;


    always @(*) begin
        
    end
endmodule