module ALU(ALU_COUT, ALUIN1, ALUIN2, ALUC);
    input ALU_COUT;

    // always @(*) begin
    // end
    
endmodule