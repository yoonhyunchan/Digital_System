module ALUcontrol(ALU_CIN, ALU_COUT);

input [4:0] ALU_CIN;
output ALU_COUT;

endmodule