module Control(ControlIn, RegWrite);


input ControlIn;
output RegWrite;

endmodule