module Shift()



endmodule