module MEM_WB ();
    
    


    always @(*) begin
        
    end
endmodule