module IF_ID();





endmodule