module SignExtended();





endmodule