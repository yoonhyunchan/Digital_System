module ALUcontrol();



endmodule