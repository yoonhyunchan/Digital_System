module ALU();
    


endmodule