module ALU(ALUIN1, ALUIN2, ALUC, ALU_OUT);
    input [31:0] ALUIN1;
    input [31:0] ALUIN2;
    input ALUC;
    output reg [31:0] ALU_OUT;


    always @(posedge ALUC) begin
    end
    
endmodule