module EX_MEM ();
    iutput reg nPC_M;
    iutput reg AOUT_M;
    iutput reg B_M;



    
endmodule