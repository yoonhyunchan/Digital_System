module tb();


endmodule