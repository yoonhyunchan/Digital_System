module and();

    input branch;
    output Zero;

    assign andout = branch & Zero;


endmodule