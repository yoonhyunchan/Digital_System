module EX_MEM ();

    input [31:0] counter1;
    input [31:0]Zero;
    input [31:0];

    output reg [31:0] nPC_M;
    output reg [31:0] AOUT_M;
    output reg [31:0] B_M;

    always @(*) begin
        
    end


endmodule