module MEM_WB ();
    
    input MDR_M;


    always @(*) begin
        
    end
endmodule