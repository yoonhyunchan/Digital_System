module SingleCpu();





endmodule