module SingleCpu(CLK, INST);
    input CLK;
    output reg INST;
    integer i;

Vr_inst_mem Vr_inst_mem1(.ADDR(ADDR), .INST(INST))







endmodule