module SignedExtension();





endmodule