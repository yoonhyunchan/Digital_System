module PC();



endmodule