module moduleName ();

reg CLK;

SingleCpu SingleCpu1 (CLK);

    
endmodule