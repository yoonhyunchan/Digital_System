module Control(ControlIn, RegWrite);




endmodule