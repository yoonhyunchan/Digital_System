module ADD_4();

    input [31:0] IN;
    output [31:0] OUT;

    assign OUT = IN +4;

endmodule