module Control(ControlIn, RegWrite);


input ControlIn;
output reg RegWrite;

endmodule