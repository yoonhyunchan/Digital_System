module tb();

    reg [11:0] input;
    wire [31:0] output;


endmodule