module ALU(ALUIN1, ALUIN2, ALUC, ALU_OUT);
    input [31:0] ALU_CIN1;
    input [31:0] ALU_CIN2;
    input ALUC;
    output reg [31:0] CLU_OUT;


    always @(posedge ALUC) begin
    end
    
endmodule