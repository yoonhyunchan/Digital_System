module ALU(ALU_COUT);
    input ALU_COUT;

    $display("%b", ALU_COUT);
endmodule