module IF_ID(Data, RST);





endmodule