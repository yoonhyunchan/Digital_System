module mux();

input ALUSrc;
input [31:0] IN1;
input [31:0] IN2;

output reg OUT;




endmodule