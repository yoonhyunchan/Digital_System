module ID_EX();


    input 


endmodule