module MEM_WB ();
    
    input [31:0] RD_mem;
    input [31:0]

    output reg [31:0] MDR_W;
    output reg [31:0] AOUT_W;


    always @(*) begin
        
    end
endmodule