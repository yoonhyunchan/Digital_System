module ALUcontrol();


endmodule