module PC();

    input [31:0] ADDR;


endmodule