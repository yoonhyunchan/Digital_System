module ALU(ALU_COUT);
    input ALU_COUT;


endmodule