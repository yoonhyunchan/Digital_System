module ALUcontrol();

input [4:0] ALU_CIN;
output ALU_COUT;

endmodule