module ALU(ALU_COUT);
    input ALU_COUT;

    // always @(*) begin
    // end
    
endmodule