module ALUcontrol();

input [4:0] ALU_CIN;

endmodule