module IF_ID(INST, Q);

    input INST;
    output reg Q;

always @(INST) begin
     Q <= INSTs;
end



endmodule