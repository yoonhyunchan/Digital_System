module EX_MEM ();
    input nPC_M;
    input AOUT_M;
    input B_M



    
endmodule