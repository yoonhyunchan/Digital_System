module SignExtended();


endmodule