module EX_MEM (
    ports
);
    
endmodule