module ALU_ADD();

input [31:0] IN1;
input [31:0] IN2;
output [31:0] Counter1;

assign 


endmodule