module tb();

    


endmodule