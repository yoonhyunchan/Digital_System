module IF_Latch();





endmodule