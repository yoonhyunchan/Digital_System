module ID_EX();

    input P_PC;
    input RD1;
    input RD2;
    input signout;



endmodule