module ID_EX();

    input P_PC;
    input RD1;
    input RD2;
    input signout;
    output P_PC2;
    output P_RD1;
    output P_RD2;
    output P_signout;


endmodule