module ALU(ALUIN1, ALUIN2, ALUC, ALU_OUT);
    input ALU_CIN;
    output reg CLU_OUT;


    always @(posedge ALUC) begin
    end
    
endmodule