module ALUcontrol(ALU_CIN, ALU_COUT);

input [3:0] ALU_CIN;
output ALU_COUT;


assign ALU_COUT = 1'b1;
endmodule